module CPU(clock, reset, 
					PCin,PCout,
					inst,
					RegWrite, ALUSrc, MemtoReg, MemRead, MemWrite, Branch,
					ALUOp,
					WriteReg,
					ReadData1, ReadData2,
					Extend64,
					ALU_B,
					ShiftOut,
					ALUCtl,
					Zero,
					ALUOut,
					AddOut,
					Add4Out,
					AndOut,
					ReadData,
					WriteData_Reg);